intent PAYMENT_INTENT
goal: "Process a payment"
inputs: "[amount: Money, account: String]"
outputs: "[id: String]"
evidence: "[legacy_code]"
tags: "[finance]"
end

mapping PAYMENT_MAPPING -> "api POST /api/payments"
request: "PaymentRequest"
response: "PaymentResponse"
end
