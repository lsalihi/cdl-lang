type Customer
  id: string
  name: string
end
